
`ifndef _tb_keydata_vh_
`define _tb_keydata_vh_

logic [31:0] KeyData1[0:612] = {
   //Start E-Matrix (100 words)      0:99  
   32'h404ecd54,      32'h719b0fa7,      32'h144fe03d,      32'h39975a62,      32'h118fdc62,     
   32'h7b6aa698,      32'h7612ab7e,      32'h038fa3c1,      32'h067ba21e,      32'h2b03703b,     
   32'h3f34b85f,      32'h558a004b,      32'h696cb6f4,      32'h5db6a195,      32'h0f4186ce,     
   32'h01146e4d,      32'h0acef1c4,      32'h32729c10,      32'h14590c6a,      32'h40e30703,     
   32'h793dd40a,      32'h663792fa,      32'h19ff6b9b,      32'h7865c658,      32'h5d85ee5a,     
   32'h2f94b11f,      32'h423462c4,      32'h0414077d,      32'h67e5617d,      32'h50f85284,     
   32'h1d89ce9c,      32'h54d90967,      32'h42a0bcf2,      32'h11fef73c,      32'h4669fb56,     
   32'h4ad00ead,      32'h7d2b228c,      32'h42f25793,      32'h1197859e,      32'h085b3260,     
   32'h18edcb23,      32'h06fa60a6,      32'h69b14b61,      32'h01eabf13,      32'h03a3bbd7,     
   32'h7269efed,      32'h2a883e68,      32'h11b0a7be,      32'h135501ae,      32'h4768f5c6,     
   32'h3fe22c29,      32'h7b5c174a,      32'h758279f2,      32'h78c70cb6,      32'h3d789ef3,     
   32'h4b25e75c,      32'h3ccda1c9,      32'h51dd7f39,      32'h0f25ff27,      32'h22c78498,     
   32'h0c2c82ff,      32'h6ddf15ce,      32'h59e1364d,      32'h5b78d25c,      32'h5e028b7b,     
   32'h5fb41263,      32'h65a765e5,      32'h3cd0350e,      32'h4f96807a,      32'h5852be38,     
   32'h02e12aae,      32'h6d17d0c8,      32'h3d0102da,      32'h6c9ddcea,      32'h34155b1e,     
   32'h6acc9fbd,      32'h4cefd3af,      32'h6324316a,      32'h04a8aca8,      32'h61d80c5b,     
   32'h7545555c,      32'h6f51fa32,      32'h78fa27a5,      32'h222b9544,      32'h113c04f6,     
   32'h7454daac,      32'h5a868c85,      32'h33963f63,      32'h524be627,      32'h73b1d9e7,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000001,     

   //Start Permutation Array (2 words) 100 : 101
   32'h00078056,      32'h00039142,     

   //Start T-Values (10 words)         102 : 111
   32'h52cfb21d,      32'h401d3c3d,      32'h06d46f6f,      32'h1b2aefd7,      32'h3080f599,     
   32'h7bf66074,      32'h3869ef5a,      32'h515e53df,      32'h72108b3d,      32'h590061d9,     

   //Start Inverse T-Values (10 words) 112 : 121
   32'h3fe2c3c2,      32'h2d304de2,      32'h0803b6b0,      32'h143f413b,      32'h71963601,     
   32'h31dd8290,      32'h1f7b0566,      32'h3bd28016,      32'h46aad12c,      32'h36c92602,     

   //Artin Generator count (1 word)  122
   32'h000008f0,   

   //Start Artin Generators, (2288 packed in 382 words)  123: 504
   32'h2b63e0e2,      32'h095b5c74,      32'h25114462,      32'h0e6b96c4,      32'h0a41ca68,     
   32'h08329226,      32'h0c735c72,      32'h226b96c5,      32'h0d29d232,      32'h265a5707,     
   32'h2d1912a4,      32'h27218c95,      32'h2d79ca34,      32'h265a1aa7,      32'h0a41c8a4,     
   32'h06288a26,      32'h24320222,      32'h24100233,      32'h2b3a4a52,      32'h07114404,     
   32'h086bd6c2,      32'h27521673,      32'h24104c54,      32'h2c8be220,      32'h0c5a1aa7,     
   32'h0648c443,      32'h0a621662,      32'h012080c7,      32'h24110c11,      32'h0c3a1464,     
   32'h2b63a295,      32'h25290474,      32'h0f6ba272,      32'h253a1ab8,      32'h0a418832,     
   32'h2c5222e6,      32'h083160e7,      32'h06210cd5,      32'h040080b4,      32'h24324833,     
   32'h020b5c01,      32'h2939ce62,      32'h02039cd5,      32'h2221c412,      32'h2642c864,     
   32'h02208005,      32'h28531d00,      32'h2b41ded5,      32'h29310401,      32'h22090674,     
   32'h26288251,      32'h00090416,      32'h2a428e41,      32'h22041f06,      32'h08210e22,     
   32'h0e5310b3,      32'h316292e6,      32'h05745f18,      32'h04300862,      32'h0541d481,     
   32'h22090673,      32'h0b208220,      32'h0a00ca64,      32'h093294d4,      32'h0b731ca4,     
   32'h06115496,      32'h2419cc54,      32'h24388220,      32'h283a90b6,      32'h227b14d7,     
   32'h26200402,      32'h066a9241,      32'h00314414,      32'h0b388041,      32'h22288e44,     
   32'h0e424653,      32'h064298e8,      32'h236b1eb4,      32'h2929c640,      32'h220b5d13,     
   32'h014ace72,      32'h24198820,      32'h08088a20,      32'h027316d6,      32'h23101072,     
   32'h02208062,      32'h0d521672,      32'h23114400,      32'h03204412,      32'h2419d053,     
   32'h00004620,      32'h07224e51,      32'h23288a20,      32'h0530c800,      32'h2d6a8021,     
   32'h04388e55,      32'h0c5b12a2,      32'h06404443,      32'h05321432,      32'h0a731274,     
   32'h241c5cc5,      32'h01194620,      32'h0008c860,      32'h23288a20,      32'h2530c811,     
   32'h27488241,      32'h22288e44,      32'h274a8640,      32'h274b56f6,      32'h2f8a9072,     
   32'h06100016,      32'h07418022,      32'h2518ce54,      32'h016ad220,      32'h24104440,     
   32'h23105693,      32'h2208c672,      32'h2d4ace92,      32'h23629a95,      32'h0118c651,     
   32'h27498032,      32'h07440442,      32'h025a5662,      32'h2249ca20,      32'h0141ca20,     
   32'h01124c51,      32'h27498432,      32'h03204402,      32'h0329d2a1,      32'h274ad8e1,     
   32'h0420c8a4,      32'h00209483,      32'h1008c871,      32'h000bdb17,      32'h0010ca64,     
   32'h253a0011,      32'h275a5ab1,      32'h0128ce54,      32'h005a56d7,      32'h00088871,     
   32'h2640c860,      32'h02200022,      32'h0221d0a1,      32'h0e108800,      32'h022192a6,     
   32'h0b7b1d00,      32'h29208864,      32'h2d524a53,      32'h2b400653,      32'h2519ca93,     
   32'h0c704400,      32'h02110c85,      32'h03324864,      32'h0c740641,      32'h0549d685,     
   32'h02190662,      32'h0113c860,      32'h26408432,      32'h0201d0a2,      32'h2f5b52a3,     
   32'h0d5a60f6,      32'h2412d262,      32'h22008493,      32'h0538c800,      32'h2d5bd874,     
   32'h02039aa4,      32'h0b498641,      32'h09390442,      32'h2c41c821,      32'h01114405,     
   32'h01829ae8,      32'h08004643,      32'h00000653,      32'h02194e85,      32'h253a54c0,     
   32'h274ad8f1,      32'h06208232,      32'h096298a4,      32'h0b41dcd5,      32'h08214c41,     
   32'h02108863,      32'h293ad2c5,      32'h01208672,      32'h074ad8f1,      32'h2d700222,     
   32'h01190e95,      32'h01194c91,      32'h2e29d0a1,      32'h2c7c52a6,      32'h10520e95,     
   32'h062c1cd7,      32'h084b98a4,      32'h04521063,      32'h06210843,      32'h02209483,     
   32'h0a418841,      32'h00018836,      32'h042084e1,      32'h08418c62,      32'h04214c43,     
   32'h04100eb4,      32'h25308a83,      32'h053a16c1,      32'h00008422,      32'h31788021,     
   32'h288bdaa6,      32'h2b499ed5,      32'h0008a0e6,      32'h2728d272,      32'h07194400,     
   32'h064a8222,      32'h25320432,      32'h29530e85,      32'h220adec7,      32'h06310402,     
   32'h07419083,      32'h047b1483,      32'h0530c823,      32'h28319ab4,      32'h24124c45,     
   32'h222a4403,      32'h2a190e80,      32'h2d710a64,      32'h285006f8,      32'h0c004653,     
   32'h293ad2d5,      32'h0a094672,      32'h007c1af8,      32'h00088871,      32'h0a08c864,     
   32'h0a60ca64,      32'h045a4eb4,      32'h02498842,      32'h22000072,      32'h2f638222,     
   32'h01629695,      32'h03298232,      32'h0549d681,      32'h27204401,      32'h2f638251,     
   32'h09101ed5,      32'h0921c443,      32'h220050b3,      32'h2328c672,      32'h09530440,     
   32'h0b7b1c43,      32'h063a90f6,      32'h033114d4,      32'h05104821,      32'h24418011,     
   32'h00000c41,      32'h0b63a041,      32'h08428c84,      32'h30735d05,      32'h06325cc5,     
   32'h2a41d8a4,      32'h02031ce8,      32'h27398a83,      32'h00090413,      32'h06404400,     
   32'h0a6990b2,      32'h0e8a98f4,      32'h0620dd16,      32'h04320422,      32'h043216c5,     
   32'h0a418821,      32'h022190a6,      32'h08110c41,      32'h0a628863,      32'h022190a6,     
   32'h022190a6,      32'h08518c22,      32'h06429843,      32'h04310422,      32'h0a6190a4,     
   32'h06410864,      32'h06429885,      32'h0e321442,      32'h0962dcd8,      32'h03315075,     
   32'h25104412,      32'h317b5693,      32'h27288000,      32'h251bdab4,      32'h251b5693,     
   32'h23395693,      32'h2d5a4e52,      32'h293ad273,      32'h2328ce51,      32'h2d5a4e51,     
   32'h235a4e51,      32'h2329d272,      32'h255a4e51,      32'h27394633,      32'h29394634,     
   32'h2518d695,      32'h2518a293,      32'h0c794633,      32'h076a92c5,      32'h0c745694,     
   32'h02200237,      32'h2c5a4e72,      32'h27294413,      32'h09304632,      32'h041a0e55,     
   32'h23104833,      32'h06414412,      32'h00110407,      32'h03298220,      32'h0c3a1453,     
   32'h2e8b1c95,      32'h2e6c1cc5,      32'h283a92c5,      32'h22090662,      32'h2b49ca51,     
   32'h2328dd16,      32'h0010ca60,      32'h28300453,      32'h27290662,      32'h2728c414,     
   32'h01110232,      32'h00198861,      32'h2a298020,      32'h28335696,      32'h262004c5,     
   32'h05104824,      32'h25208011,      32'h22288252,      32'h24104c43,      32'h0642c620,     
   32'h0d42cc82,      32'h08310415,      32'h00000c42,      32'h0d838820,      32'h00110c85,     
   32'h09508a74,      32'h0a6c6043,      32'h262ad064,      32'h2749ca41,      32'h2b49ca52,     
   32'h275b62f6,      32'h29395ab4,      32'h254ad295,      32'h25394620,      32'h2b49ca31,     
   32'h293ad2f6,      32'h29395ab4,      32'h0d5a5694,      32'h09194eb5,      32'h064a92c5,     
   32'h0e7a1672,      32'h0620cc06,      32'h04326022,      32'h047a1673,      32'h04320443,     
   32'h0e834401,      32'h272190a6,      32'h0809d0a6,      32'h04300441,      32'h08531d01,     
   32'h2c500443,      32'h2a6a1464,      32'h03399262,      32'h04300440,      32'h064298e1,     
   32'h08530022,      32'h08590443,      32'h012190a6,      32'h06008a81,      32'h08531c02,     
   32'h0b800443,      32'h09208864,      32'h04195683,      32'h24390693,      32'h08500441,     
   32'h01390443,      32'h085b9a51,      32'h08538ec3,      32'h0f6298e3,      32'h0a3262f6,     
   32'h283b5496,      32'h000002d5,        

   
   //SHA 256 Hash bytes (8 words)  
   32'h72e97ea4,      32'h5e7103d5,      32'hd09e3350,      32'hcc58e359,      32'h11e9191c,      
   32'haea36116,      32'h9adb036e,      32'h41976058,     

   //Public Matrix prime (100 words)  
   32'h170d63b4,      32'h233802cd,      32'h137fbb9f,      32'h2e2d9a3d,      32'h18e96ff7,     
   32'h0c88294d,      32'h42f95e19,      32'h05eeb23b,      32'h5d7cc700,      32'h5c4c4f7c,     
   32'h3be98ddd,      32'h6785f9c2,      32'h048592b6,      32'h19102992,      32'h4186d083,     
   32'h34d76d36,      32'h25eeac32,      32'h65cc812e,      32'h195b5590,      32'h269d1ec9,     
   32'h4a169d6c,      32'h7d2473f6,      32'h3824df2c,      32'h60c69eb6,      32'h0906ca9c,     
   32'h780d24b7,      32'h1858ef53,      32'h56d2d406,      32'h311d6c0b,      32'h0c5cdc10,     
   32'h1e42fb6c,      32'h6d2dd2c0,      32'h562db687,      32'h6c9c885d,      32'h734f8dd5,     
   32'h78e7c06b,      32'h5bc31a10,      32'h7683518f,      32'h67e2ef83,      32'h1809452d,     
   32'h7a7eb3de,      32'h2425210f,      32'h5fd3dc2a,      32'h6bcde8fb,      32'h7bf5c5ae,     
   32'h055901d8,      32'h072571c7,      32'h3f600d47,      32'h13ebf95e,      32'h49c8c99b,     
   32'h479b5a39,      32'h409d5de9,      32'h49b2132d,      32'h43879cb3,      32'h52941e33,     
   32'h0dbd6407,      32'h4f6ec4ad,      32'h10da38f3,      32'h27bb3af7,      32'h3d927d94,     
   32'h16296f72,      32'h6ee4bf58,      32'h6dddeba7,      32'h610ab329,      32'h36086709,     
   32'h1156e1c2,      32'h26cd6af4,      32'h7dea5e8f,      32'h24897681,      32'h233a3c75,     
   32'h375998f5,      32'h51a078ed,      32'h2b503db5,      32'h4cfe7432,      32'h44d6360b,     
   32'h2f5e7ffb,      32'h1c7461bb,      32'h1ec5f288,      32'h4e6a40ef,      32'h54463191,     
   32'h2b6aeccf,      32'h1e7d9d92,      32'h1dac8962,      32'h2247c64b,      32'h3e3f793b,     
   32'h55a0207d,      32'h5caacc61,      32'h1e749fa8,      32'h3fdee368,      32'h36c2b686,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000001     
  
};


logic [31:0] SIGNATURE[0:504] = {

   //Start E-Matrix (100 words)        
   32'h404ecd54,      32'h719b0fa7,      32'h144fe03d,      32'h39975a62,      32'h118fdc62,     
   32'h7b6aa698,      32'h7612ab7e,      32'h038fa3c1,      32'h067ba21e,      32'h2b03703b,     
   32'h3f34b85f,      32'h558a004b,      32'h696cb6f4,      32'h5db6a195,      32'h0f4186ce,     
   32'h01146e4d,      32'h0acef1c4,      32'h32729c10,      32'h14590c6a,      32'h40e30703,     
   32'h793dd40a,      32'h663792fa,      32'h19ff6b9b,      32'h7865c658,      32'h5d85ee5a,     
   32'h2f94b11f,      32'h423462c4,      32'h0414077d,      32'h67e5617d,      32'h50f85284,     
   32'h1d89ce9c,      32'h54d90967,      32'h42a0bcf2,      32'h11fef73c,      32'h4669fb56,     
   32'h4ad00ead,      32'h7d2b228c,      32'h42f25793,      32'h1197859e,      32'h085b3260,     
   32'h18edcb23,      32'h06fa60a6,      32'h69b14b61,      32'h01eabf13,      32'h03a3bbd7,     
   32'h7269efed,      32'h2a883e68,      32'h11b0a7be,      32'h135501ae,      32'h4768f5c6,     
   32'h3fe22c29,      32'h7b5c174a,      32'h758279f2,      32'h78c70cb6,      32'h3d789ef3,     
   32'h4b25e75c,      32'h3ccda1c9,      32'h51dd7f39,      32'h0f25ff27,      32'h22c78498,     
   32'h0c2c82ff,      32'h6ddf15ce,      32'h59e1364d,      32'h5b78d25c,      32'h5e028b7b,     
   32'h5fb41263,      32'h65a765e5,      32'h3cd0350e,      32'h4f96807a,      32'h5852be38,     
   32'h02e12aae,      32'h6d17d0c8,      32'h3d0102da,      32'h6c9ddcea,      32'h34155b1e,     
   32'h6acc9fbd,      32'h4cefd3af,      32'h6324316a,      32'h04a8aca8,      32'h61d80c5b,     
   32'h7545555c,      32'h6f51fa32,      32'h78fa27a5,      32'h222b9544,      32'h113c04f6,     
   32'h7454daac,      32'h5a868c85,      32'h33963f63,      32'h524be627,      32'h73b1d9e7,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000001,     

   //Start Permutation Array (2 words) 
   32'h00078056,      32'h00039142,     

   //Start T-Values (10 words)         
   32'h52cfb21d,      32'h401d3c3d,      32'h06d46f6f,      32'h1b2aefd7,      32'h3080f599,     
   32'h7bf66074,      32'h3869ef5a,      32'h515e53df,      32'h72108b3d,      32'h590061d9,     

   //Start Inverse T-Values (10 words) 
   32'h3fe2c3c2,      32'h2d304de2,      32'h0803b6b0,      32'h143f413b,      32'h71963601,     
   32'h31dd8290,      32'h1f7b0566,      32'h3bd28016,      32'h46aad12c,      32'h36c92602,     

   //Artin Generator count (1 word)  
   32'h000008f0,   

   //Start Artin Generators, (2288 packed in 382 words) 
   32'h2b63e0e2,      32'h095b5c74,      32'h25114462,      32'h0e6b96c4,      32'h0a41ca68,     
   32'h08329226,      32'h0c735c72,      32'h226b96c5,      32'h0d29d232,      32'h265a5707,     
   32'h2d1912a4,      32'h27218c95,      32'h2d79ca34,      32'h265a1aa7,      32'h0a41c8a4,     
   32'h06288a26,      32'h24320222,      32'h24100233,      32'h2b3a4a52,      32'h07114404,     
   32'h086bd6c2,      32'h27521673,      32'h24104c54,      32'h2c8be220,      32'h0c5a1aa7,     
   32'h0648c443,      32'h0a621662,      32'h012080c7,      32'h24110c11,      32'h0c3a1464,     
   32'h2b63a295,      32'h25290474,      32'h0f6ba272,      32'h253a1ab8,      32'h0a418832,     
   32'h2c5222e6,      32'h083160e7,      32'h06210cd5,      32'h040080b4,      32'h24324833,     
   32'h020b5c01,      32'h2939ce62,      32'h02039cd5,      32'h2221c412,      32'h2642c864,     
   32'h02208005,      32'h28531d00,      32'h2b41ded5,      32'h29310401,      32'h22090674,     
   32'h26288251,      32'h00090416,      32'h2a428e41,      32'h22041f06,      32'h08210e22,     
   32'h0e5310b3,      32'h316292e6,      32'h05745f18,      32'h04300862,      32'h0541d481,     
   32'h22090673,      32'h0b208220,      32'h0a00ca64,      32'h093294d4,      32'h0b731ca4,     
   32'h06115496,      32'h2419cc54,      32'h24388220,      32'h283a90b6,      32'h227b14d7,     
   32'h26200402,      32'h066a9241,      32'h00314414,      32'h0b388041,      32'h22288e44,     
   32'h0e424653,      32'h064298e8,      32'h236b1eb4,      32'h2929c640,      32'h220b5d13,     
   32'h014ace72,      32'h24198820,      32'h08088a20,      32'h027316d6,      32'h23101072,     
   32'h02208062,      32'h0d521672,      32'h23114400,      32'h03204412,      32'h2419d053,     
   32'h00004620,      32'h07224e51,      32'h23288a20,      32'h0530c800,      32'h2d6a8021,     
   32'h04388e55,      32'h0c5b12a2,      32'h06404443,      32'h05321432,      32'h0a731274,     
   32'h241c5cc5,      32'h01194620,      32'h0008c860,      32'h23288a20,      32'h2530c811,     
   32'h27488241,      32'h22288e44,      32'h274a8640,      32'h274b56f6,      32'h2f8a9072,     
   32'h06100016,      32'h07418022,      32'h2518ce54,      32'h016ad220,      32'h24104440,     
   32'h23105693,      32'h2208c672,      32'h2d4ace92,      32'h23629a95,      32'h0118c651,     
   32'h27498032,      32'h07440442,      32'h025a5662,      32'h2249ca20,      32'h0141ca20,     
   32'h01124c51,      32'h27498432,      32'h03204402,      32'h0329d2a1,      32'h274ad8e1,     
   32'h0420c8a4,      32'h00209483,      32'h1008c871,      32'h000bdb17,      32'h0010ca64,     
   32'h253a0011,      32'h275a5ab1,      32'h0128ce54,      32'h005a56d7,      32'h00088871,     
   32'h2640c860,      32'h02200022,      32'h0221d0a1,      32'h0e108800,      32'h022192a6,     
   32'h0b7b1d00,      32'h29208864,      32'h2d524a53,      32'h2b400653,      32'h2519ca93,     
   32'h0c704400,      32'h02110c85,      32'h03324864,      32'h0c740641,      32'h0549d685,     
   32'h02190662,      32'h0113c860,      32'h26408432,      32'h0201d0a2,      32'h2f5b52a3,     
   32'h0d5a60f6,      32'h2412d262,      32'h22008493,      32'h0538c800,      32'h2d5bd874,     
   32'h02039aa4,      32'h0b498641,      32'h09390442,      32'h2c41c821,      32'h01114405,     
   32'h01829ae8,      32'h08004643,      32'h00000653,      32'h02194e85,      32'h253a54c0,     
   32'h274ad8f1,      32'h06208232,      32'h096298a4,      32'h0b41dcd5,      32'h08214c41,     
   32'h02108863,      32'h293ad2c5,      32'h01208672,      32'h074ad8f1,      32'h2d700222,     
   32'h01190e95,      32'h01194c91,      32'h2e29d0a1,      32'h2c7c52a6,      32'h10520e95,     
   32'h062c1cd7,      32'h084b98a4,      32'h04521063,      32'h06210843,      32'h02209483,     
   32'h0a418841,      32'h00018836,      32'h042084e1,      32'h08418c62,      32'h04214c43,     
   32'h04100eb4,      32'h25308a83,      32'h053a16c1,      32'h00008422,      32'h31788021,     
   32'h288bdaa6,      32'h2b499ed5,      32'h0008a0e6,      32'h2728d272,      32'h07194400,     
   32'h064a8222,      32'h25320432,      32'h29530e85,      32'h220adec7,      32'h06310402,     
   32'h07419083,      32'h047b1483,      32'h0530c823,      32'h28319ab4,      32'h24124c45,     
   32'h222a4403,      32'h2a190e80,      32'h2d710a64,      32'h285006f8,      32'h0c004653,     
   32'h293ad2d5,      32'h0a094672,      32'h007c1af8,      32'h00088871,      32'h0a08c864,     
   32'h0a60ca64,      32'h045a4eb4,      32'h02498842,      32'h22000072,      32'h2f638222,     
   32'h01629695,      32'h03298232,      32'h0549d681,      32'h27204401,      32'h2f638251,     
   32'h09101ed5,      32'h0921c443,      32'h220050b3,      32'h2328c672,      32'h09530440,     
   32'h0b7b1c43,      32'h063a90f6,      32'h033114d4,      32'h05104821,      32'h24418011,     
   32'h00000c41,      32'h0b63a041,      32'h08428c84,      32'h30735d05,      32'h06325cc5,     
   32'h2a41d8a4,      32'h02031ce8,      32'h27398a83,      32'h00090413,      32'h06404400,     
   32'h0a6990b2,      32'h0e8a98f4,      32'h0620dd16,      32'h04320422,      32'h043216c5,     
   32'h0a418821,      32'h022190a6,      32'h08110c41,      32'h0a628863,      32'h022190a6,     
   32'h022190a6,      32'h08518c22,      32'h06429843,      32'h04310422,      32'h0a6190a4,     
   32'h06410864,      32'h06429885,      32'h0e321442,      32'h0962dcd8,      32'h03315075,     
   32'h25104412,      32'h317b5693,      32'h27288000,      32'h251bdab4,      32'h251b5693,     
   32'h23395693,      32'h2d5a4e52,      32'h293ad273,      32'h2328ce51,      32'h2d5a4e51,     
   32'h235a4e51,      32'h2329d272,      32'h255a4e51,      32'h27394633,      32'h29394634,     
   32'h2518d695,      32'h2518a293,      32'h0c794633,      32'h076a92c5,      32'h0c745694,     
   32'h02200237,      32'h2c5a4e72,      32'h27294413,      32'h09304632,      32'h041a0e55,     
   32'h23104833,      32'h06414412,      32'h00110407,      32'h03298220,      32'h0c3a1453,     
   32'h2e8b1c95,      32'h2e6c1cc5,      32'h283a92c5,      32'h22090662,      32'h2b49ca51,     
   32'h2328dd16,      32'h0010ca60,      32'h28300453,      32'h27290662,      32'h2728c414,     
   32'h01110232,      32'h00198861,      32'h2a298020,      32'h28335696,      32'h262004c5,     
   32'h05104824,      32'h25208011,      32'h22288252,      32'h24104c43,      32'h0642c620,     
   32'h0d42cc82,      32'h08310415,      32'h00000c42,      32'h0d838820,      32'h00110c85,     
   32'h09508a74,      32'h0a6c6043,      32'h262ad064,      32'h2749ca41,      32'h2b49ca52,     
   32'h275b62f6,      32'h29395ab4,      32'h254ad295,      32'h25394620,      32'h2b49ca31,     
   32'h293ad2f6,      32'h29395ab4,      32'h0d5a5694,      32'h09194eb5,      32'h064a92c5,     
   32'h0e7a1672,      32'h0620cc06,      32'h04326022,      32'h047a1673,      32'h04320443,     
   32'h0e834401,      32'h272190a6,      32'h0809d0a6,      32'h04300441,      32'h08531d01,     
   32'h2c500443,      32'h2a6a1464,      32'h03399262,      32'h04300440,      32'h064298e1,     
   32'h08530022,      32'h08590443,      32'h012190a6,      32'h06008a81,      32'h08531c02,     
   32'h0b800443,      32'h09208864,      32'h04195683,      32'h24390693,      32'h08500441,     
   32'h01390443,      32'h085b9a51,      32'h08538ec3,      32'h0f6298e3,      32'h0a3262f6,     
   32'h283b5496,      32'h000002d5        
};


logic [31:0] ENCODER[0:204] = {

   //Start E-Matrix (100 words)        
   32'h00000001,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000001,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000001,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000001,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000001,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000001,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000001,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000001,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000001,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,     
   32'h00000000,      32'h00000000,      32'h00000000,      32'h00000000,      32'h00000001,     

   //Start Permutation Array (2 words) 
   32'h00043210,      32'h00098765,     

   //Start T-Values (10 words)         
   32'h52cfb21d,      32'h401d3c3d,      32'h06d46f6f,      32'h1b2aefd7,      32'h3080f599,     
   32'h7bf66074,      32'h3869ef5a,      32'h515e53df,      32'h72108b3d,      32'h590061d9,     

   //Start Inverse T-Values (10 words) 
   32'h3fe2c3c2,      32'h2d304de2,      32'h0803b6b0,      32'h143f413b,      32'h71963601,     
   32'h31dd8290,      32'h1f7b0566,      32'h3bd28016,      32'h46aad12c,      32'h36c92602,     

   //Artin Generator count (1 word)  
   32'h000001ea,   

   //Start Artin Generators, (490 packed in 82 words) 
   32'h084298e8,      32'h0a639ed5,      32'h00008864,      32'h2c5a4e51,      32'h0a63a117,     
   32'h064210a5,      32'h0e7b5483,      32'h0c5298c6,      32'h064294a6,      32'h24108842,     
   32'h28319093,      32'h0a5298d5,      32'h0e7b5484,      32'h022190a6,      32'h06394400,     
   32'h02108842,      32'h29394400,      32'h0e841ed5,      32'h063190a6,      32'h2d5a0c42,     
   32'h0a63a117,      32'h02218c64,      32'h29390400,      32'h064298d5,      32'h0a635683,     
   32'h042190a5,      32'h0e7b5693,      32'h022190a6,      32'h29394400,      32'h0a639ed5,     
   32'h06319084,      32'h24100022,      32'h117b5693,      32'h064298e8,      32'h29390422,     
   32'h064298d5,      32'h09390422,      32'h06420c64,      32'h29390422,      32'h0e845ed5,     
   32'h064294a6,      32'h25100022,      32'h0e7b5693,      32'h064210a6,      32'h06319083,     
   32'h02218c42,      32'h28394400,      32'h0e845ed5,      32'h084294a6,      32'h04218c64,     
   32'h06319083,      32'h0d5a0c42,      32'h022190a6,      32'h0d5a4e41,      32'h0a6314a6,     
   32'h0a5298c5,      32'h00008864,      32'h2d5a4e51,      32'h084298e7,      32'h022190a5,     
   32'h06394400,      32'h04218c42,      32'h0a631693,      32'h2c520c64,      32'h0a63a117,     
   32'h2d520c64,      32'h064298e7,      32'h02108842,      32'h29394400,      32'h0a639ed5,     
   32'h0a631484,      32'h064210a5,      32'h00008422,      32'h0d5a0e51,      32'h063190a6,     
   32'h2d5a4c42,      32'h084298e7,      32'h022190a5,      32'h09390400,      32'h06420c64,     
   32'h29390422,      32'h000c5ed5        
};


`endif
